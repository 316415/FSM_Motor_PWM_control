`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/10/14 13:00:40
// Design Name: 
// Module Name: FND_2x4_decoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module FND_position_decoder(
    input i_clk,
    output o_position
    );

    reg r_position = 1'b0;
    assign o_position = r_position;
endmodule
